`default_nettype none
module instrconunit(
   input Clock,
   input Reset,
   input BRANCH,
   input JUMP,
   input [7:0] imm,
   output [7:0] PC
);

endmodule
