`default_nettype none
module Hardware(
   input CLK,
   input RST,
   input [3:0] H,
   output [3:0] V,
   output [3:0] SD,
   output [7:0] SEG,
   output [7:0] LD,
   input [7:0] SB,
   output Buzz
`ifdef SIMULATION
   ,
   output [7:0] io_ena,
   inout [7:0] io_0,
   inout [7:0] io_1,
   inout [7:0] io_2,
   inout [7:0] io_3,
   inout [7:0] io_4,
   inout [7:0] io_5,
   inout [7:0] io_6,
   inout [7:0] io_7
`endif
   );

   // fundamental modules
   wire Clock, Reset;
   assign Clock = CLK;
   rst_recover rst(Clock, RST, Reset);

   // links
   wire [7:0] ou_L, ou_H;
`ifndef SIMULATION
   wire [7:0] io_ena;
   wire [7:0] io_0, io_1, io_2, io_3;
   wire [7:0] io_4, io_5, io_6, io_7;
`endif

   // auxillary
   latch_buffer lat0(
      .Clock(Clock), .Reset(Reset),
      .en(io_ena[0]), .in(io_0), .out(ou_L));
   latch_buffer lat1(
      .Clock(Clock), .Reset(Reset),
      .en(io_ena[1]), .in(io_1), .out(ou_H));
   latch_buffer lat7(
      .Clock(Clock), .Reset(Reset),
      .en(io_ena[7]), .in(io_7), .out(LD));

   assign Buzz = ~LD[0];

   // main modules
   CPU u(
      .Clock(Clock), .Reset(Reset),
      .io_ena(io_ena),
      .io_0(io_0), .io_1(io_1),
      .io_2(io_2), .io_3(io_3),
      .io_4(io_4), .io_5(io_5),
      .io_6(io_6), .io_7(io_7));

   Input in(
      .Clock(Clock), .Reset(Reset),
      .H(H), .V(V), .ack(io_ena[2]),
      .io(io_2));

   seg out(
      .CLK_seg(Clock),
      .data_inH(ou_H), .data_inL(ou_L),
      .seg_sel(SD), .data_out(SEG));

endmodule
