`default_nettype none
module lpm_rom_256_16(
   input Clock,
   input Reset,
   input [7:0] address,
   output [15:0] q
);

endmodule
