`default_nettype none
module ctrlunit(
   input [3:0] OP,
   input ZERO,
   output JUMP,
   output BRANCH,
   output [2:0] ALUC,
   output ALUSRCB,
   output WRITEMEM,
   output WRITEREG,
   output MEMTOREG,
   output REGDES,
   output WRFLAG
);

endmodule
