`default_nettype none
module Flag(
   input Clock,
   input Reset,
   input [7:0] Flagin,
   output [7:0] Flagout
);

endmodule
